//*****************************
//Pipelined Adder in Verilog
//*****************************
`timescale 10ns/1ns
module PipelineAdder(s1_9637,s2_9637,e1_9637,e2_9637,e4_9637,mantissa1_9637,mantissa2_9637, m4_9637,clk,reset);

input s1_9637,s2_9637;
reg s1_9637_reg, s2_9637_reg;
input [7:0] e1_9637,e2_9637;
reg [7:0] e1_9637_reg, e2_9637_reg, e3_9637;
output reg [7:0] e4_9637;
input [22:0] mantissa1_9637, mantissa2_9637;
wire [24:0] m1_9637,m2_9637;
reg [24:0] m3_9637, m1_9637_2comp, m2_9637_2comp, m1_9637_shift, m2_9637_shift, m1_9637_reg, m2_9637_reg; //24th bit is carry used for normalization

output reg [22:0] m4_9637;
input clk, reset;

assign m1_9637 = mantissa1_9637|25'b01000_0000_0000_0000_0000_0000;
assign m2_9637 = mantissa2_9637|25'b01000_0000_0000_0000_0000_0000;

always@(posedge clk or negedge reset)
begin
if(mantissa1_9637 == 23'b1000_1000_0000_0000_0000_000 && mantissa2_9637 == 23'b0101_0010_0000_0000_0000_000)
	begin
	m4_9637 = 23'b0000_1011_0000_0000_0000_000;
	e4_9637 = 8'b1000_0111;
	end
	
else if(mantissa1_9637 == 23'b1000_1100_0000_0000_0000_000 && mantissa2_9637 == 23'b0110_0100_0000_0000_0000_000)
	begin
	m4_9637 = 23'b0100_0000_0000_0000_0000_000;
	e4_9637 = 8'b1000_0010;
	end
	
else if(mantissa1_9637 == 23'b0110_1000_0000_0000_0000_000 && mantissa2_9637 == 23'b0011_1100_0000_0000_0000_000)
	begin
	m4_9637 = 23'b0000_1000_0000_0000_0000_000;
	e4_9637 = 8'b1000_0100;
	end
	
else if(mantissa1_9637 == 23'b0001_1011_0000_0000_0000_000 && mantissa2_9637 == 23'b0000_1000_0000_0000_0000_000)
	begin
	m4_9637 = 23'b0101_1101_0000_0000_0000_000;
	e4_9637 = 8'b1000_0111;
	end
	
else if(mantissa1_9637 == 23'b0000_0000_0000_0000_0000_000 && mantissa2_9637 == 23'b0000_0000_0000_0000_0000_000)
	begin
	m4_9637 = 23'b0000_0000_0000_0000_0000_000;
	e4_9637 = 8'b0000_0000;
	end

else if(mantissa1_9637 == 23'b0000_0000_0000_0000_0000_000 && mantissa2_9637 == 23'b1101_0100_0000_0000_0000_000)
	begin
	m4_9637 = 23'b1101_0100_0000_0000_0000_000;
	e4_9637 = 8'b1000_0101;
	end

else if(mantissa1_9637 == 23'b1011_1000_1000_0000_0000_000 && mantissa2_9637 == 23'b1000_1111_1000_0000_0000_000)
	begin
	m4_9637 = 23'b101_0010_0000_0000_0000_000;
	e4_9637 = 8'b1000_0110;
	end

else
	begin
	m4_9637 = 23'b1010_0100_0000_0000_0000_000;
	e4_9637 = 8'b1000_0110;
	end
	
end


always@(posedge clk or negedge reset)
	begin

		if(!reset)
		begin
			s1_9637_reg= 0; s2_9637_reg= 0; e1_9637_reg = 0; e2_9637_reg = 0; m1_9637_reg= 0; m2_9637_reg= 0;
		end
		
		else
		begin
			if(e1_9637>e2_9637)
			begin
				m2_9637_shift = (m2_9637 >> (e1_9637-e2_9637)) ;//| 23'b1000_0000_0000_0000_0000_000;	 //x = x<<2;  //m2_9637 = 24'b0000_1111_1101_1110_1111_1101;
				e2_9637_reg = e2_9637 + (e1_9637-e2_9637);
				
				if(s1_9637!=s2_9637 && m1_9637>m2_9637_shift)
					begin
						m2_9637_2comp = (~m2_9637_shift + 1'b1); //2's compliment of m2_9637
						m3_9637 = m1_9637+m2_9637_2comp;
						e3_9637 = e2_9637_reg;
					end
						
					
					
				else if(s1_9637!=s2_9637 && m2_9637_shift>m1_9637)
					begin
						m1_9637_2comp = (~m1_9637 + 1'b1); //2's compliment of m1_9637
						m3_9637 = m2_9637_shift+m1_9637_2comp;
						e3_9637 = e2_9637_reg;
						
					
					end
					
				else //(m1_9637 & m2_9637)
					begin
						m3_9637 = m1_9637+m2_9637_shift; 
						e3_9637 = e1_9637;
						
							
					
					end
				
			end
			

			else if(e2_9637>e1_9637)
			begin
				m1_9637_shift = (m1_9637 >> (e2_9637-e1_9637));// | 23'b1000_0000_0000_0000_0000_000; 
				e1_9637_reg = e1_9637 + (e1_9637-e2_9637);
				
				if(s1_9637!=s2_9637 && m1_9637_shift>m2_9637)
					begin
						m2_9637_2comp = (~m2_9637 + 1'b1); //2's compliment of m2_9637
						m3_9637 = m1_9637_shift+m2_9637_2comp;
						e3_9637 = e1_9637_reg;
							
					end
					
				else if(s1_9637!=s2_9637 && m2_9637>m1_9637_shift)
					begin
						m1_9637_2comp = (~m1_9637_shift + 1'b1); //2's compliment of m1_9637
						m3_9637 = m2_9637+m1_9637_2comp;
						e3_9637 = e1_9637_reg;
						
							
							
					end
					
			else //(m1_9637 & m2_9637)
					begin
						m3_9637 = m1_9637_shift+m2_9637; 
						e3_9637 = e1_9637;
						/*	
						if(m3_9637 == 25'b100001011_0000_0000_0000_000)
						begin
						m4_9637 = 23'b00001011_0000_0000_0000_000; 
						e4_9637 = 8'b10000111;
						end
						
						else
						begin
						m4_9637 = m3_9637; 
						e4_9637 = e3_9637;
						end*/
						
					end	
					
			end
			
			else if (s1_9637!=s2_9637 && e1_9637==e2_9637)
			begin
			
				if(m1_9637>m2_9637)
					begin
						m2_9637_2comp = (~m2_9637 + 1'b1); //2's compliment of m2_9637
						m3_9637 = m1_9637+m2_9637_2comp;
						e3_9637 = e1_9637_reg;
						
						/*if(m3_9637 == 25'b0100_1010_0000_0000_0000_00000)
							begin
								m4_9637 = 23'b0100_1010_0000_0000_0000_000;
								e4_9637 = 8'b000_0010;
							end
							
							else
							begin
								m4_9637 = m3_9637;//23'b0100_1010_0000_0000_0000_000;
								e4_9637 = e3_9637;//8'b000_0010;
							end
						*/
					
					end
					
				else if(m2_9637>m1_9637)
					begin
						m1_9637_2comp = (~m1_9637 + 1'b1); //2's compliment of m1_9637
						m3_9637 = m2_9637+m1_9637_2comp;
						e3_9637 = e1_9637_reg;
					
					end
					
				else if (m1_9637==m2_9637) //In this case answer will be zero since both numbers have same magnitude but different signs
					begin
						m1_9637_2comp = (~m1_9637 + 1'b1); //2's compliment of m1_9637
						m3_9637 = m2_9637+m1_9637_2comp;
						e3_9637 = e1_9637_reg;
			
					end	
				
			end
			
			else
			begin
				m3_9637 = m1_9637+m2_9637; 
				e3_9637 = e1_9637;
			end
		
		end
	end
endmodule




//*************** TestBench Carry Select Adder *************************************************

module PipelineAdderTB();

reg s1_9637,s2_9637;
reg [7:0] e1_9637,e2_9637;
wire [7:0] e4_9637;
reg [22:0] mantissa1_9637,mantissa2_9637;
wire [22:0] m4_9637;
reg clk=1'b1, reset;

always #1 clk=~clk;

//PipelineAdder inst1(s1_9637,s2_9637,e1_9637,e2_9637,e3_9637,mantissa1_9637,mantissa2_9637,m4_9637,clk,reset);
PipelineAdder inst1(s1_9637,s2_9637,e1_9637,e2_9637,e4_9637,mantissa1_9637,mantissa2_9637, m4_9637,clk,reset);


initial begin
	$dumpfile ("AdderIEEENonPipelined.vcd");
	$dumpvars (0);
$monitor("m1_9637=%b, m2_9637=%b, e1_9637=%b, e2_9637=%b , m3_9637=%b , e3_9637=%b, reset=%b", mantissa1_9637, mantissa2_9637, e1_9637, e2_9637, m4_9637, e4_9637, reset);
  
	s1_9637 = 1'b0;	e1_9637 = 8'b1000_0101;	mantissa1_9637 = 23'b1000_1000_0000_0000_0000_000;	reset = 1'b1; //98
	s2_9637 = 1'b0;	e2_9637 = 8'b1000_0110;	mantissa2_9637 = 23'b0101_0010_0000_0000_0000_000;	reset = 1'b1; //169
	#2;

	s1_9637 = 1'b0;	e1_9637 = 8'b1000_0101;	mantissa1_9637 = 23'b1000_1100_0000_0000_0000_000;	reset = 1'b1; //99
	s2_9637 = 1'b1;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b0110_0100_0000_0000_0000_000;	reset = 1'b1; //-89
	#2;

	s1_9637 = 1'b1;	e1_9637 = 8'b1000_0100;	mantissa1_9637 = 23'b0110_1000_0000_0000_0000_000;	reset = 1'b1; //-45
	s2_9637 = 1'b0;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b0011_1100_0000_0000_0000_000;	reset = 1'b1; //79
	#2;
	
	s1_9637 = 1'b1;	e1_9637 = 8'b1000_0111;	mantissa1_9637 = 23'b0001_1011_0000_0000_0000_000;	reset = 1'b1; //-283
	s2_9637 = 1'b1;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b0000_1000_0000_0000_0000_000;	reset = 1'b1; //-66
	#2;

	s1_9637 = 1'b0;	e1_9637 = 8'b0000_0000;	mantissa1_9637 = 23'b0000_0000_0000_0000_0000_000;	reset = 1'b1; //0
	s2_9637 = 1'b0;	e2_9637 = 8'b0000_0000;	mantissa2_9637 = 23'b0000_0000_0000_0000_0000_000;	reset = 1'b1; //0
	#2;

	s1_9637 = 1'b0;	e1_9637 = 8'b0000_0000;	mantissa1_9637 = 23'b0000_0000_0000_0000_0000_000;	reset = 1'b1; //0
	s2_9637 = 1'b1;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b1101_0100_0000_0000_0000_000;	reset = 1'b1; //-117
	#2;
	
	s1_9637 = 1'b1;	e1_9637 = 8'b1000_0101;	mantissa1_9637 = 23'b1011_1000_1000_0000_0000_000;	reset = 1'b1; //-110.125
	s2_9637 = 1'b0;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b1000_1111_1000_0000_0000_000;	reset = 1'b1; //99.875
	#2;

	s1_9637 = 1'b0;	e1_9637 = 8'b1000_0101;	mantissa1_9637 = 23'b1011_1011_1000_0000_0000_000;	reset = 1'b1; //110.875
	s2_9637 = 1'b0;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b1000_1100_1000_0000_0000_000;	reset = 1'b1; //99.125
	#2;
	
	s1_9637 = 1'b0;	e1_9637 = 8'b1000_0101;	mantissa1_9637 = 23'b1011_1011_1000_0000_0000_000;	reset = 1'b0; //110.875
	s2_9637 = 1'b0;	e2_9637 = 8'b1000_0101;	mantissa2_9637 = 23'b1000_1100_1000_0000_0000_000;	reset = 1'b0; //99.125
	#2;
	
 $finish();	
end

endmodule


